library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_unsigned.ALL;

entity l_conv is
	Port (clk : in STD_LOGIC;
	load : in STD_LOGIC; 
	dinL : in STD_LOGIC_VECTOR (127 downto 0); 
	fin_outL : out STD_LOGIC_VECTOR (127 downto 0);
	fin_out_stbL : out STD_LOGIC );
end l_conv;

architecture Behavioral of l_conv is
    type Tmem is array (0 to 255) of std_logic_vector(7 downto 0);
    constant FG148: Tmem:= (0 => x"00", 1 => x"94", 2 => x"eb", 3 => x"7f", 4 => x"15", 5 => x"81", 6 => x"fe", 7 => x"6a", 8 => x"2a", 9 => x"be", 10 => x"c1", 11 => x"55", 12 => x"3f", 13 => x"ab", 14 => x"d4", 15 => x"40", 16 => x"54", 17 => x"c0", 18 => x"bf", 19 => x"2b", 20 => x"41", 21 => x"d5", 22 => x"aa", 23 => x"3e", 24 => x"7e", 25 => x"ea", 26 => x"95", 27 => x"01", 28 => x"6b", 29 => x"ff", 30 => x"80", 31 => x"14", 32 => x"a8", 33 => x"3c", 34 => x"43", 35 => x"d7", 36 => x"bd", 37 => x"29", 38 => x"56", 39 => x"c2", 40 => x"82", 41 => x"16", 42 => x"69", 43 => x"fd", 44 => x"97", 45 => x"03", 46 => x"7c", 47 => x"e8", 48 => x"fc", 49 => x"68", 50 => x"17", 51 => x"83", 52 => x"e9", 53 => x"7d", 54 => x"02", 55 => x"96", 56 => x"d6", 57 => x"42", 58 => x"3d", 59 => x"a9", 60 => x"c3", 61 => x"57", 62 => x"28", 63 => x"bc", 64 => x"93", 65 => x"07", 66 => x"78", 67 => x"ec", 68 => x"86", 69 => x"12", 70 => x"6d", 71 => x"f9", 72 => x"b9", 73 => x"2d", 74 => x"52", 75 => x"c6", 76 => x"ac", 77 => x"38", 78 => x"47", 79 => x"d3", 80 => x"c7", 81 => x"53", 82 => x"2c", 83 => x"b8", 84 => x"d2", 85 => x"46", 86 => x"39", 87 => x"ad", 88 => x"ed", 89 => x"79", 90 => x"06", 91 => x"92", 92 => x"f8", 93 => x"6c", 94 => x"13", 95 => x"87", 96 => x"3b", 97 => x"af", 98 => x"d0", 99 => x"44", 100 => x"2e", 101 => x"ba", 102 => x"c5", 103 => x"51", 104 => x"11", 105 => x"85", 106 => x"fa", 107 => x"6e", 108 => x"04", 109 => x"90", 110 => x"ef", 111 => x"7b", 112 => x"6f", 113 => x"fb", 114 => x"84", 115 => x"10", 116 => x"7a", 117 => x"ee", 118 => x"91", 119 => x"05", 120 => x"45", 121 => x"d1", 122 => x"ae", 123 => x"3a", 124 => x"50", 125 => x"c4", 126 => x"bb", 127 => x"2f", 128 => x"e5", 129 => x"71", 130 => x"0e", 131 => x"9a", 132 => x"f0", 133 => x"64", 134 => x"1b", 135 => x"8f", 136 => x"cf", 137 => x"5b", 138 => x"24", 139 => x"b0", 140 => x"da", 141 => x"4e", 142 => x"31", 143 => x"a5", 144 => x"b1", 145 => x"25", 146 => x"5a", 147 => x"ce", 148 => x"a4", 149 => x"30", 150 => x"4f", 151 => x"db", 152 => x"9b", 153 => x"0f", 154 => x"70", 155 => x"e4", 156 => x"8e", 157 => x"1a", 158 => x"65", 159 => x"f1", 160 => x"4d", 161 => x"d9", 162 => x"a6", 163 => x"32", 164 => x"58", 165 => x"cc", 166 => x"b3", 167 => x"27", 168 => x"67", 169 => x"f3", 170 => x"8c", 171 => x"18", 172 => x"72", 173 => x"e6", 174 => x"99", 175 => x"0d", 176 => x"19", 177 => x"8d", 178 => x"f2", 179 => x"66", 180 => x"0c", 181 => x"98", 182 => x"e7", 183 => x"73", 184 => x"33", 185 => x"a7", 186 => x"d8", 187 => x"4c", 188 => x"26", 189 => x"b2", 190 => x"cd", 191 => x"59", 192 => x"76", 193 => x"e2", 194 => x"9d", 195 => x"09", 196 => x"63", 197 => x"f7", 198 => x"88", 199 => x"1c", 200 => x"5c", 201 => x"c8", 202 => x"b7", 203 => x"23", 204 => x"49", 205 => x"dd", 206 => x"a2", 207 => x"36", 208 => x"22", 209 => x"b6", 210 => x"c9", 211 => x"5d", 212 => x"37", 213 => x"a3", 214 => x"dc", 215 => x"48", 216 => x"08", 217 => x"9c", 218 => x"e3", 219 => x"77", 220 => x"1d", 221 => x"89", 222 => x"f6", 223 => x"62", 224 => x"de", 225 => x"4a", 226 => x"35", 227 => x"a1", 228 => x"cb", 229 => x"5f", 230 => x"20", 231 => x"b4", 232 => x"f4", 233 => x"60", 234 => x"1f", 235 => x"8b", 236 => x"e1", 237 => x"75", 238 => x"0a", 239 => x"9e", 240 => x"8a", 241 => x"1e", 242 => x"61", 243 => x"f5", 244 => x"9f", 245 => x"0b", 246 => x"74", 247 => x"e0", 248 => x"a0", 249 => x"34", 250 => x"4b", 251 => x"df", 252 => x"b5", 253 => x"21", 254 => x"5e", 255 => x"ca");
    constant FG32: Tmem:= (0 => x"00", 1 => x"20", 2 => x"40", 3 => x"60", 4 => x"80", 5 => x"a0", 6 => x"c0", 7 => x"e0", 8 => x"c3", 9 => x"e3", 10 => x"83", 11 => x"a3", 12 => x"43", 13 => x"63", 14 => x"03", 15 => x"23", 16 => x"45", 17 => x"65", 18 => x"05", 19 => x"25", 20 => x"c5", 21 => x"e5", 22 => x"85", 23 => x"a5", 24 => x"86", 25 => x"a6", 26 => x"c6", 27 => x"e6", 28 => x"06", 29 => x"26", 30 => x"46", 31 => x"66", 32 => x"8a", 33 => x"aa", 34 => x"ca", 35 => x"ea", 36 => x"0a", 37 => x"2a", 38 => x"4a", 39 => x"6a", 40 => x"49", 41 => x"69", 42 => x"09", 43 => x"29", 44 => x"c9", 45 => x"e9", 46 => x"89", 47 => x"a9", 48 => x"cf", 49 => x"ef", 50 => x"8f", 51 => x"af", 52 => x"4f", 53 => x"6f", 54 => x"0f", 55 => x"2f", 56 => x"0c", 57 => x"2c", 58 => x"4c", 59 => x"6c", 60 => x"8c", 61 => x"ac", 62 => x"cc", 63 => x"ec", 64 => x"d7", 65 => x"f7", 66 => x"97", 67 => x"b7", 68 => x"57", 69 => x"77", 70 => x"17", 71 => x"37", 72 => x"14", 73 => x"34", 74 => x"54", 75 => x"74", 76 => x"94", 77 => x"b4", 78 => x"d4", 79 => x"f4", 80 => x"92", 81 => x"b2", 82 => x"d2", 83 => x"f2", 84 => x"12", 85 => x"32", 86 => x"52", 87 => x"72", 88 => x"51", 89 => x"71", 90 => x"11", 91 => x"31", 92 => x"d1", 93 => x"f1", 94 => x"91", 95 => x"b1", 96 => x"5d", 97 => x"7d", 98 => x"1d", 99 => x"3d", 100 => x"dd", 101 => x"fd", 102 => x"9d", 103 => x"bd", 104 => x"9e", 105 => x"be", 106 => x"de", 107 => x"fe", 108 => x"1e", 109 => x"3e", 110 => x"5e", 111 => x"7e", 112 => x"18", 113 => x"38", 114 => x"58", 115 => x"78", 116 => x"98", 117 => x"b8", 118 => x"d8", 119 => x"f8", 120 => x"db", 121 => x"fb", 122 => x"9b", 123 => x"bb", 124 => x"5b", 125 => x"7b", 126 => x"1b", 127 => x"3b", 128 => x"6d", 129 => x"4d", 130 => x"2d", 131 => x"0d", 132 => x"ed", 133 => x"cd", 134 => x"ad", 135 => x"8d", 136 => x"ae", 137 => x"8e", 138 => x"ee", 139 => x"ce", 140 => x"2e", 141 => x"0e", 142 => x"6e", 143 => x"4e", 144 => x"28", 145 => x"08", 146 => x"68", 147 => x"48", 148 => x"a8", 149 => x"88", 150 => x"e8", 151 => x"c8", 152 => x"eb", 153 => x"cb", 154 => x"ab", 155 => x"8b", 156 => x"6b", 157 => x"4b", 158 => x"2b", 159 => x"0b", 160 => x"e7", 161 => x"c7", 162 => x"a7", 163 => x"87", 164 => x"67", 165 => x"47", 166 => x"27", 167 => x"07", 168 => x"24", 169 => x"04", 170 => x"64", 171 => x"44", 172 => x"a4", 173 => x"84", 174 => x"e4", 175 => x"c4", 176 => x"a2", 177 => x"82", 178 => x"e2", 179 => x"c2", 180 => x"22", 181 => x"02", 182 => x"62", 183 => x"42", 184 => x"61", 185 => x"41", 186 => x"21", 187 => x"01", 188 => x"e1", 189 => x"c1", 190 => x"a1", 191 => x"81", 192 => x"ba", 193 => x"9a", 194 => x"fa", 195 => x"da", 196 => x"3a", 197 => x"1a", 198 => x"7a", 199 => x"5a", 200 => x"79", 201 => x"59", 202 => x"39", 203 => x"19", 204 => x"f9", 205 => x"d9", 206 => x"b9", 207 => x"99", 208 => x"ff", 209 => x"df", 210 => x"bf", 211 => x"9f", 212 => x"7f", 213 => x"5f", 214 => x"3f", 215 => x"1f", 216 => x"3c", 217 => x"1c", 218 => x"7c", 219 => x"5c", 220 => x"bc", 221 => x"9c", 222 => x"fc", 223 => x"dc", 224 => x"30", 225 => x"10", 226 => x"70", 227 => x"50", 228 => x"b0", 229 => x"90", 230 => x"f0", 231 => x"d0", 232 => x"f3", 233 => x"d3", 234 => x"b3", 235 => x"93", 236 => x"73", 237 => x"53", 238 => x"33", 239 => x"13", 240 => x"75", 241 => x"55", 242 => x"35", 243 => x"15", 244 => x"f5", 245 => x"d5", 246 => x"b5", 247 => x"95", 248 => x"b6", 249 => x"96", 250 => x"f6", 251 => x"d6", 252 => x"36", 253 => x"16", 254 => x"76", 255 => x"56");
    constant FG133: Tmem:= (0 => x"00", 1 => x"85", 2 => x"c9", 3 => x"4c", 4 => x"51", 5 => x"d4", 6 => x"98", 7 => x"1d", 8 => x"a2", 9 => x"27", 10 => x"6b", 11 => x"ee", 12 => x"f3", 13 => x"76", 14 => x"3a", 15 => x"bf", 16 => x"87", 17 => x"02", 18 => x"4e", 19 => x"cb", 20 => x"d6", 21 => x"53", 22 => x"1f", 23 => x"9a", 24 => x"25", 25 => x"a0", 26 => x"ec", 27 => x"69", 28 => x"74", 29 => x"f1", 30 => x"bd", 31 => x"38", 32 => x"cd", 33 => x"48", 34 => x"04", 35 => x"81", 36 => x"9c", 37 => x"19", 38 => x"55", 39 => x"d0", 40 => x"6f", 41 => x"ea", 42 => x"a6", 43 => x"23", 44 => x"3e", 45 => x"bb", 46 => x"f7", 47 => x"72", 48 => x"4a", 49 => x"cf", 50 => x"83", 51 => x"06", 52 => x"1b", 53 => x"9e", 54 => x"d2", 55 => x"57", 56 => x"e8", 57 => x"6d", 58 => x"21", 59 => x"a4", 60 => x"b9", 61 => x"3c", 62 => x"70", 63 => x"f5", 64 => x"59", 65 => x"dc", 66 => x"90", 67 => x"15", 68 => x"08", 69 => x"8d", 70 => x"c1", 71 => x"44", 72 => x"fb", 73 => x"7e", 74 => x"32", 75 => x"b7", 76 => x"aa", 77 => x"2f", 78 => x"63", 79 => x"e6", 80 => x"de", 81 => x"5b", 82 => x"17", 83 => x"92", 84 => x"8f", 85 => x"0a", 86 => x"46", 87 => x"c3", 88 => x"7c", 89 => x"f9", 90 => x"b5", 91 => x"30", 92 => x"2d", 93 => x"a8", 94 => x"e4", 95 => x"61", 96 => x"94", 97 => x"11", 98 => x"5d", 99 => x"d8", 100 => x"c5", 101 => x"40", 102 => x"0c", 103 => x"89", 104 => x"36", 105 => x"b3", 106 => x"ff", 107 => x"7a", 108 => x"67", 109 => x"e2", 110 => x"ae", 111 => x"2b", 112 => x"13", 113 => x"96", 114 => x"da", 115 => x"5f", 116 => x"42", 117 => x"c7", 118 => x"8b", 119 => x"0e", 120 => x"b1", 121 => x"34", 122 => x"78", 123 => x"fd", 124 => x"e0", 125 => x"65", 126 => x"29", 127 => x"ac", 128 => x"b2", 129 => x"37", 130 => x"7b", 131 => x"fe", 132 => x"e3", 133 => x"66", 134 => x"2a", 135 => x"af", 136 => x"10", 137 => x"95", 138 => x"d9", 139 => x"5c", 140 => x"41", 141 => x"c4", 142 => x"88", 143 => x"0d", 144 => x"35", 145 => x"b0", 146 => x"fc", 147 => x"79", 148 => x"64", 149 => x"e1", 150 => x"ad", 151 => x"28", 152 => x"97", 153 => x"12", 154 => x"5e", 155 => x"db", 156 => x"c6", 157 => x"43", 158 => x"0f", 159 => x"8a", 160 => x"7f", 161 => x"fa", 162 => x"b6", 163 => x"33", 164 => x"2e", 165 => x"ab", 166 => x"e7", 167 => x"62", 168 => x"dd", 169 => x"58", 170 => x"14", 171 => x"91", 172 => x"8c", 173 => x"09", 174 => x"45", 175 => x"c0", 176 => x"f8", 177 => x"7d", 178 => x"31", 179 => x"b4", 180 => x"a9", 181 => x"2c", 182 => x"60", 183 => x"e5", 184 => x"5a", 185 => x"df", 186 => x"93", 187 => x"16", 188 => x"0b", 189 => x"8e", 190 => x"c2", 191 => x"47", 192 => x"eb", 193 => x"6e", 194 => x"22", 195 => x"a7", 196 => x"ba", 197 => x"3f", 198 => x"73", 199 => x"f6", 200 => x"49", 201 => x"cc", 202 => x"80", 203 => x"05", 204 => x"18", 205 => x"9d", 206 => x"d1", 207 => x"54", 208 => x"6c", 209 => x"e9", 210 => x"a5", 211 => x"20", 212 => x"3d", 213 => x"b8", 214 => x"f4", 215 => x"71", 216 => x"ce", 217 => x"4b", 218 => x"07", 219 => x"82", 220 => x"9f", 221 => x"1a", 222 => x"56", 223 => x"d3", 224 => x"26", 225 => x"a3", 226 => x"ef", 227 => x"6a", 228 => x"77", 229 => x"f2", 230 => x"be", 231 => x"3b", 232 => x"84", 233 => x"01", 234 => x"4d", 235 => x"c8", 236 => x"d5", 237 => x"50", 238 => x"1c", 239 => x"99", 240 => x"a1", 241 => x"24", 242 => x"68", 243 => x"ed", 244 => x"f0", 245 => x"75", 246 => x"39", 247 => x"bc", 248 => x"03", 249 => x"86", 250 => x"ca", 251 => x"4f", 252 => x"52", 253 => x"d7", 254 => x"9b", 255 => x"1e");
    constant FG16: Tmem:= (0 => x"00", 1 => x"10", 2 => x"20", 3 => x"30", 4 => x"40", 5 => x"50", 6 => x"60", 7 => x"70", 8 => x"80", 9 => x"90", 10 => x"a0", 11 => x"b0", 12 => x"c0", 13 => x"d0", 14 => x"e0", 15 => x"f0", 16 => x"c3", 17 => x"d3", 18 => x"e3", 19 => x"f3", 20 => x"83", 21 => x"93", 22 => x"a3", 23 => x"b3", 24 => x"43", 25 => x"53", 26 => x"63", 27 => x"73", 28 => x"03", 29 => x"13", 30 => x"23", 31 => x"33", 32 => x"45", 33 => x"55", 34 => x"65", 35 => x"75", 36 => x"05", 37 => x"15", 38 => x"25", 39 => x"35", 40 => x"c5", 41 => x"d5", 42 => x"e5", 43 => x"f5", 44 => x"85", 45 => x"95", 46 => x"a5", 47 => x"b5", 48 => x"86", 49 => x"96", 50 => x"a6", 51 => x"b6", 52 => x"c6", 53 => x"d6", 54 => x"e6", 55 => x"f6", 56 => x"06", 57 => x"16", 58 => x"26", 59 => x"36", 60 => x"46", 61 => x"56", 62 => x"66", 63 => x"76", 64 => x"8a", 65 => x"9a", 66 => x"aa", 67 => x"ba", 68 => x"ca", 69 => x"da", 70 => x"ea", 71 => x"fa", 72 => x"0a", 73 => x"1a", 74 => x"2a", 75 => x"3a", 76 => x"4a", 77 => x"5a", 78 => x"6a", 79 => x"7a", 80 => x"49", 81 => x"59", 82 => x"69", 83 => x"79", 84 => x"09", 85 => x"19", 86 => x"29", 87 => x"39", 88 => x"c9", 89 => x"d9", 90 => x"e9", 91 => x"f9", 92 => x"89", 93 => x"99", 94 => x"a9", 95 => x"b9", 96 => x"cf", 97 => x"df", 98 => x"ef", 99 => x"ff", 100 => x"8f", 101 => x"9f", 102 => x"af", 103 => x"bf", 104 => x"4f", 105 => x"5f", 106 => x"6f", 107 => x"7f", 108 => x"0f", 109 => x"1f", 110 => x"2f", 111 => x"3f", 112 => x"0c", 113 => x"1c", 114 => x"2c", 115 => x"3c", 116 => x"4c", 117 => x"5c", 118 => x"6c", 119 => x"7c", 120 => x"8c", 121 => x"9c", 122 => x"ac", 123 => x"bc", 124 => x"cc", 125 => x"dc", 126 => x"ec", 127 => x"fc", 128 => x"d7", 129 => x"c7", 130 => x"f7", 131 => x"e7", 132 => x"97", 133 => x"87", 134 => x"b7", 135 => x"a7", 136 => x"57", 137 => x"47", 138 => x"77", 139 => x"67", 140 => x"17", 141 => x"07", 142 => x"37", 143 => x"27", 144 => x"14", 145 => x"04", 146 => x"34", 147 => x"24", 148 => x"54", 149 => x"44", 150 => x"74", 151 => x"64", 152 => x"94", 153 => x"84", 154 => x"b4", 155 => x"a4", 156 => x"d4", 157 => x"c4", 158 => x"f4", 159 => x"e4", 160 => x"92", 161 => x"82", 162 => x"b2", 163 => x"a2", 164 => x"d2", 165 => x"c2", 166 => x"f2", 167 => x"e2", 168 => x"12", 169 => x"02", 170 => x"32", 171 => x"22", 172 => x"52", 173 => x"42", 174 => x"72", 175 => x"62", 176 => x"51", 177 => x"41", 178 => x"71", 179 => x"61", 180 => x"11", 181 => x"01", 182 => x"31", 183 => x"21", 184 => x"d1", 185 => x"c1", 186 => x"f1", 187 => x"e1", 188 => x"91", 189 => x"81", 190 => x"b1", 191 => x"a1", 192 => x"5d", 193 => x"4d", 194 => x"7d", 195 => x"6d", 196 => x"1d", 197 => x"0d", 198 => x"3d", 199 => x"2d", 200 => x"dd", 201 => x"cd", 202 => x"fd", 203 => x"ed", 204 => x"9d", 205 => x"8d", 206 => x"bd", 207 => x"ad", 208 => x"9e", 209 => x"8e", 210 => x"be", 211 => x"ae", 212 => x"de", 213 => x"ce", 214 => x"fe", 215 => x"ee", 216 => x"1e", 217 => x"0e", 218 => x"3e", 219 => x"2e", 220 => x"5e", 221 => x"4e", 222 => x"7e", 223 => x"6e", 224 => x"18", 225 => x"08", 226 => x"38", 227 => x"28", 228 => x"58", 229 => x"48", 230 => x"78", 231 => x"68", 232 => x"98", 233 => x"88", 234 => x"b8", 235 => x"a8", 236 => x"d8", 237 => x"c8", 238 => x"f8", 239 => x"e8", 240 => x"db", 241 => x"cb", 242 => x"fb", 243 => x"eb", 244 => x"9b", 245 => x"8b", 246 => x"bb", 247 => x"ab", 248 => x"5b", 249 => x"4b", 250 => x"7b", 251 => x"6b", 252 => x"1b", 253 => x"0b", 254 => x"3b", 255 => x"2b");
    constant FG194: Tmem:= (0 => x"00", 1 => x"c2", 2 => x"47", 3 => x"85", 4 => x"8e", 5 => x"4c", 6 => x"c9", 7 => x"0b", 8 => x"df", 9 => x"1d", 10 => x"98", 11 => x"5a", 12 => x"51", 13 => x"93", 14 => x"16", 15 => x"d4", 16 => x"7d", 17 => x"bf", 18 => x"3a", 19 => x"f8", 20 => x"f3", 21 => x"31", 22 => x"b4", 23 => x"76", 24 => x"a2", 25 => x"60", 26 => x"e5", 27 => x"27", 28 => x"2c", 29 => x"ee", 30 => x"6b", 31 => x"a9", 32 => x"fa", 33 => x"38", 34 => x"bd", 35 => x"7f", 36 => x"74", 37 => x"b6", 38 => x"33", 39 => x"f1", 40 => x"25", 41 => x"e7", 42 => x"62", 43 => x"a0", 44 => x"ab", 45 => x"69", 46 => x"ec", 47 => x"2e", 48 => x"87", 49 => x"45", 50 => x"c0", 51 => x"02", 52 => x"09", 53 => x"cb", 54 => x"4e", 55 => x"8c", 56 => x"58", 57 => x"9a", 58 => x"1f", 59 => x"dd", 60 => x"d6", 61 => x"14", 62 => x"91", 63 => x"53", 64 => x"37", 65 => x"f5", 66 => x"70", 67 => x"b2", 68 => x"b9", 69 => x"7b", 70 => x"fe", 71 => x"3c", 72 => x"e8", 73 => x"2a", 74 => x"af", 75 => x"6d", 76 => x"66", 77 => x"a4", 78 => x"21", 79 => x"e3", 80 => x"4a", 81 => x"88", 82 => x"0d", 83 => x"cf", 84 => x"c4", 85 => x"06", 86 => x"83", 87 => x"41", 88 => x"95", 89 => x"57", 90 => x"d2", 91 => x"10", 92 => x"1b", 93 => x"d9", 94 => x"5c", 95 => x"9e", 96 => x"cd", 97 => x"0f", 98 => x"8a", 99 => x"48", 100 => x"43", 101 => x"81", 102 => x"04", 103 => x"c6", 104 => x"12", 105 => x"d0", 106 => x"55", 107 => x"97", 108 => x"9c", 109 => x"5e", 110 => x"db", 111 => x"19", 112 => x"b0", 113 => x"72", 114 => x"f7", 115 => x"35", 116 => x"3e", 117 => x"fc", 118 => x"79", 119 => x"bb", 120 => x"6f", 121 => x"ad", 122 => x"28", 123 => x"ea", 124 => x"e1", 125 => x"23", 126 => x"a6", 127 => x"64", 128 => x"6e", 129 => x"ac", 130 => x"29", 131 => x"eb", 132 => x"e0", 133 => x"22", 134 => x"a7", 135 => x"65", 136 => x"b1", 137 => x"73", 138 => x"f6", 139 => x"34", 140 => x"3f", 141 => x"fd", 142 => x"78", 143 => x"ba", 144 => x"13", 145 => x"d1", 146 => x"54", 147 => x"96", 148 => x"9d", 149 => x"5f", 150 => x"da", 151 => x"18", 152 => x"cc", 153 => x"0e", 154 => x"8b", 155 => x"49", 156 => x"42", 157 => x"80", 158 => x"05", 159 => x"c7", 160 => x"94", 161 => x"56", 162 => x"d3", 163 => x"11", 164 => x"1a", 165 => x"d8", 166 => x"5d", 167 => x"9f", 168 => x"4b", 169 => x"89", 170 => x"0c", 171 => x"ce", 172 => x"c5", 173 => x"07", 174 => x"82", 175 => x"40", 176 => x"e9", 177 => x"2b", 178 => x"ae", 179 => x"6c", 180 => x"67", 181 => x"a5", 182 => x"20", 183 => x"e2", 184 => x"36", 185 => x"f4", 186 => x"71", 187 => x"b3", 188 => x"b8", 189 => x"7a", 190 => x"ff", 191 => x"3d", 192 => x"59", 193 => x"9b", 194 => x"1e", 195 => x"dc", 196 => x"d7", 197 => x"15", 198 => x"90", 199 => x"52", 200 => x"86", 201 => x"44", 202 => x"c1", 203 => x"03", 204 => x"08", 205 => x"ca", 206 => x"4f", 207 => x"8d", 208 => x"24", 209 => x"e6", 210 => x"63", 211 => x"a1", 212 => x"aa", 213 => x"68", 214 => x"ed", 215 => x"2f", 216 => x"fb", 217 => x"39", 218 => x"bc", 219 => x"7e", 220 => x"75", 221 => x"b7", 222 => x"32", 223 => x"f0", 224 => x"a3", 225 => x"61", 226 => x"e4", 227 => x"26", 228 => x"2d", 229 => x"ef", 230 => x"6a", 231 => x"a8", 232 => x"7c", 233 => x"be", 234 => x"3b", 235 => x"f9", 236 => x"f2", 237 => x"30", 238 => x"b5", 239 => x"77", 240 => x"de", 241 => x"1c", 242 => x"99", 243 => x"5b", 244 => x"50", 245 => x"92", 246 => x"17", 247 => x"d5", 248 => x"01", 249 => x"c3", 250 => x"46", 251 => x"84", 252 => x"8f", 253 => x"4d", 254 => x"c8", 255 => x"0a");
    constant FG192: Tmem:= ( 0 => x"00", 1 => x"c0", 2 => x"43", 3 => x"83", 4 => x"86", 5 => x"46", 6 => x"c5", 7 => x"05", 8 => x"cf", 9 => x"0f", 10 => x"8c", 11 => x"4c", 12 => x"49", 13 => x"89", 14 => x"0a", 15 => x"ca", 16 => x"5d", 17 => x"9d", 18 => x"1e", 19 => x"de", 20 => x"db", 21 => x"1b", 22 => x"98", 23 => x"58", 24 => x"92", 25 => x"52", 26 => x"d1", 27 => x"11", 28 => x"14", 29 => x"d4", 30 => x"57", 31 => x"97", 32 => x"ba", 33 => x"7a", 34 => x"f9", 35 => x"39", 36 => x"3c", 37 => x"fc", 38 => x"7f", 39 => x"bf", 40 => x"75", 41 => x"b5", 42 => x"36", 43 => x"f6", 44 => x"f3", 45 => x"33", 46 => x"b0", 47 => x"70", 48 => x"e7", 49 => x"27", 50 => x"a4", 51 => x"64", 52 => x"61", 53 => x"a1", 54 => x"22", 55 => x"e2", 56 => x"28", 57 => x"e8", 58 => x"6b", 59 => x"ab", 60 => x"ae", 61 => x"6e", 62 => x"ed", 63 => x"2d", 64 => x"b7", 65 => x"77", 66 => x"f4", 67 => x"34", 68 => x"31", 69 => x"f1", 70 => x"72", 71 => x"b2", 72 => x"78", 73 => x"b8", 74 => x"3b", 75 => x"fb", 76 => x"fe", 77 => x"3e", 78 => x"bd", 79 => x"7d", 80 => x"ea", 81 => x"2a", 82 => x"a9", 83 => x"69", 84 => x"6c", 85 => x"ac", 86 => x"2f", 87 => x"ef", 88 => x"25", 89 => x"e5", 90 => x"66", 91 => x"a6", 92 => x"a3", 93 => x"63", 94 => x"e0", 95 => x"20", 96 => x"0d", 97 => x"cd", 98 => x"4e", 99 => x"8e", 100 => x"8b", 101 => x"4b", 102 => x"c8", 103 => x"08", 104 => x"c2", 105 => x"02", 106 => x"81", 107 => x"41", 108 => x"44", 109 => x"84", 110 => x"07", 111 => x"c7", 112 => x"50", 113 => x"90", 114 => x"13", 115 => x"d3", 116 => x"d6", 117 => x"16", 118 => x"95", 119 => x"55", 120 => x"9f", 121 => x"5f", 122 => x"dc", 123 => x"1c", 124 => x"19", 125 => x"d9", 126 => x"5a", 127 => x"9a", 128 => x"ad", 129 => x"6d", 130 => x"ee", 131 => x"2e", 132 => x"2b", 133 => x"eb", 134 => x"68", 135 => x"a8", 136 => x"62", 137 => x"a2", 138 => x"21", 139 => x"e1", 140 => x"e4", 141 => x"24", 142 => x"a7", 143 => x"67", 144 => x"f0", 145 => x"30", 146 => x"b3", 147 => x"73", 148 => x"76", 149 => x"b6", 150 => x"35", 151 => x"f5", 152 => x"3f", 153 => x"ff", 154 => x"7c", 155 => x"bc", 156 => x"b9", 157 => x"79", 158 => x"fa", 159 => x"3a", 160 => x"17", 161 => x"d7", 162 => x"54", 163 => x"94", 164 => x"91", 165 => x"51", 166 => x"d2", 167 => x"12", 168 => x"d8", 169 => x"18", 170 => x"9b", 171 => x"5b", 172 => x"5e", 173 => x"9e", 174 => x"1d", 175 => x"dd", 176 => x"4a", 177 => x"8a", 178 => x"09", 179 => x"c9", 180 => x"cc", 181 => x"0c", 182 => x"8f", 183 => x"4f", 184 => x"85", 185 => x"45", 186 => x"c6", 187 => x"06", 188 => x"03", 189 => x"c3", 190 => x"40", 191 => x"80", 192 => x"1a", 193 => x"da", 194 => x"59", 195 => x"99", 196 => x"9c", 197 => x"5c", 198 => x"df", 199 => x"1f", 200 => x"d5", 201 => x"15", 202 => x"96", 203 => x"56", 204 => x"53", 205 => x"93", 206 => x"10", 207 => x"d0", 208 => x"47", 209 => x"87", 210 => x"04", 211 => x"c4", 212 => x"c1", 213 => x"01", 214 => x"82", 215 => x"42", 216 => x"88", 217 => x"48", 218 => x"cb", 219 => x"0b", 220 => x"0e", 221 => x"ce", 222 => x"4d", 223 => x"8d", 224 => x"a0", 225 => x"60", 226 => x"e3", 227 => x"23", 228 => x"26", 229 => x"e6", 230 => x"65", 231 => x"a5", 232 => x"6f", 233 => x"af", 234 => x"2c", 235 => x"ec", 236 => x"e9", 237 => x"29", 238 => x"aa", 239 => x"6a", 240 => x"fd", 241 => x"3d", 242 => x"be", 243 => x"7e", 244 => x"7b", 245 => x"bb", 246 => x"38", 247 => x"f8", 248 => x"32", 249 => x"f2", 250 => x"71", 251 => x"b1", 252 => x"b4", 253 => x"74", 254 => x"f7", 255 => x"37");
    constant FG251: Tmem:= ( 0 => x"00", 1 => x"fb", 2 => x"35", 3 => x"ce", 4 => x"6a", 5 => x"91", 6 => x"5f", 7 => x"a4", 8 => x"d4", 9 => x"2f", 10 => x"e1", 11 => x"1a", 12 => x"be", 13 => x"45", 14 => x"8b", 15 => x"70", 16 => x"6b", 17 => x"90", 18 => x"5e", 19 => x"a5", 20 => x"01", 21 => x"fa", 22 => x"34", 23 => x"cf", 24 => x"bf", 25 => x"44", 26 => x"8a", 27 => x"71", 28 => x"d5", 29 => x"2e", 30 => x"e0", 31 => x"1b", 32 => x"d6", 33 => x"2d", 34 => x"e3", 35 => x"18", 36 => x"bc", 37 => x"47", 38 => x"89", 39 => x"72", 40 => x"02", 41 => x"f9", 42 => x"37", 43 => x"cc", 44 => x"68", 45 => x"93", 46 => x"5d", 47 => x"a6", 48 => x"bd", 49 => x"46", 50 => x"88", 51 => x"73", 52 => x"d7", 53 => x"2c", 54 => x"e2", 55 => x"19", 56 => x"69", 57 => x"92", 58 => x"5c", 59 => x"a7", 60 => x"03", 61 => x"f8", 62 => x"36", 63 => x"cd", 64 => x"6f", 65 => x"94", 66 => x"5a", 67 => x"a1", 68 => x"05", 69 => x"fe", 70 => x"30", 71 => x"cb", 72 => x"bb", 73 => x"40", 74 => x"8e", 75 => x"75", 76 => x"d1", 77 => x"2a", 78 => x"e4", 79 => x"1f", 80 => x"04", 81 => x"ff", 82 => x"31", 83 => x"ca", 84 => x"6e", 85 => x"95", 86 => x"5b", 87 => x"a0", 88 => x"d0", 89 => x"2b", 90 => x"e5", 91 => x"1e", 92 => x"ba", 93 => x"41", 94 => x"8f", 95 => x"74", 96 => x"b9", 97 => x"42", 98 => x"8c", 99 => x"77", 100 => x"d3", 101 => x"28", 102 => x"e6", 103 => x"1d", 104 => x"6d", 105 => x"96", 106 => x"58", 107 => x"a3", 108 => x"07", 109 => x"fc", 110 => x"32", 111 => x"c9", 112 => x"d2", 113 => x"29", 114 => x"e7", 115 => x"1c", 116 => x"b8", 117 => x"43", 118 => x"8d", 119 => x"76", 120 => x"06", 121 => x"fd", 122 => x"33", 123 => x"c8", 124 => x"6c", 125 => x"97", 126 => x"59", 127 => x"a2", 128 => x"de", 129 => x"25", 130 => x"eb", 131 => x"10", 132 => x"b4", 133 => x"4f", 134 => x"81", 135 => x"7a", 136 => x"0a", 137 => x"f1", 138 => x"3f", 139 => x"c4", 140 => x"60", 141 => x"9b", 142 => x"55", 143 => x"ae", 144 => x"b5", 145 => x"4e", 146 => x"80", 147 => x"7b", 148 => x"df", 149 => x"24", 150 => x"ea", 151 => x"11", 152 => x"61", 153 => x"9a", 154 => x"54", 155 => x"af", 156 => x"0b", 157 => x"f0", 158 => x"3e", 159 => x"c5", 160 => x"08", 161 => x"f3", 162 => x"3d", 163 => x"c6", 164 => x"62", 165 => x"99", 166 => x"57", 167 => x"ac", 168 => x"dc", 169 => x"27", 170 => x"e9", 171 => x"12", 172 => x"b6", 173 => x"4d", 174 => x"83", 175 => x"78", 176 => x"63", 177 => x"98", 178 => x"56", 179 => x"ad", 180 => x"09", 181 => x"f2", 182 => x"3c", 183 => x"c7", 184 => x"b7", 185 => x"4c", 186 => x"82", 187 => x"79", 188 => x"dd", 189 => x"26", 190 => x"e8", 191 => x"13", 192 => x"b1", 193 => x"4a", 194 => x"84", 195 => x"7f", 196 => x"db", 197 => x"20", 198 => x"ee", 199 => x"15", 200 => x"65", 201 => x"9e", 202 => x"50", 203 => x"ab", 204 => x"0f", 205 => x"f4", 206 => x"3a", 207 => x"c1", 208 => x"da", 209 => x"21", 210 => x"ef", 211 => x"14", 212 => x"b0", 213 => x"4b", 214 => x"85", 215 => x"7e", 216 => x"0e", 217 => x"f5", 218 => x"3b", 219 => x"c0", 220 => x"64", 221 => x"9f", 222 => x"51", 223 => x"aa", 224 => x"67", 225 => x"9c", 226 => x"52", 227 => x"a9", 228 => x"0d", 229 => x"f6", 230 => x"38", 231 => x"c3", 232 => x"b3", 233 => x"48", 234 => x"86", 235 => x"7d", 236 => x"d9", 237 => x"22", 238 => x"ec", 239 => x"17", 240 => x"0c", 241 => x"f7", 242 => x"39", 243 => x"c2", 244 => x"66", 245 => x"9d", 246 => x"53", 247 => x"a8", 248 => x"d8", 249 => x"23", 250 => x"ed", 251 => x"16", 252 => x"b2", 253 => x"49", 254 => x"87", 255 => x"7c");
	signal tmpL: std_logic_vector(127 downto 0) := (others => '0');
	signal countL: std_logic_vector(4 downto 0) := "00000";
	signal work: std_logic := '0';
	
begin
process(clk)
variable i0, i1, i2, i3, i4, i5, i7, i9, i10, i11, i12, i13, i14 : integer;
begin
if (clk'event and clk ='1') then
	if (load = '1') then
		tmpL<=dinL;
		countL <= "00000";
		work <= '1';
		fin_out_stbL <= '0';
	else
		if(countL(4) = '0' ) then
			fin_out_stbL <= '0';
			if (work = '1') then
			i0 := CONV_INTEGER(tmpL(119 downto 112));
			i1 := CONV_INTEGER(tmpL(111 downto 104));
			i2 := CONV_INTEGER(tmpL(103 downto 96));
			i3 := CONV_INTEGER(tmpL(95 downto 88));
			i4 := CONV_INTEGER(tmpL(87 downto 80));
			i5 := CONV_INTEGER(tmpL(79 downto 72));
			
			i7 := CONV_INTEGER(tmpL(63 downto 56));
			
			i9 := CONV_INTEGER(tmpL(47 downto 40));
			i10 := CONV_INTEGER(tmpL(39 downto 32));
			i11 := CONV_INTEGER(tmpL(31 downto 24));
			i12 := CONV_INTEGER(tmpL(23 downto 16));
			i13 := CONV_INTEGER(tmpL(15 downto 8));
			i14 := CONV_INTEGER(tmpL(7 downto 0));
			
			tmpL <=  tmpL(119 downto 0) & (FG148(i0) xor FG32(i1) xor FG133(i2) xor FG16(i3) xor FG194(i4) xor FG192(i5) xor tmpL(71 downto 64) xor FG251(i7) xor tmpL(55 downto 48) xor FG192(i9) xor FG194(i10) xor FG16(i11) xor FG133(i12) xor FG32(i13) xor FG148(i14) xor tmpL(127 downto 120)) ;
			countL <= countL + 1;
			end if;
		else
			fin_out_stbL <= '1';
			countL <= "00000";
			work <= '0';
		end if;
	end if;
end if;
end process;
fin_outL <= tmpL;
end Behavioral;